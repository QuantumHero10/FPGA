module lts1 (
    input [7:0] SW,
	 output [7:0] LED
);
    assign LED = SW;
endmodule
