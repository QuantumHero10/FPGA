`timescale 1ns/1ns

module muon(
input wire clk,
input wire reset,
input wire signal,
input wire [5:0] switch,
output wire [7:0] led,
output wire [7:0] gpio,
output wire [5:0] gpiob,
output wire [7:0] count
);

reg [9:0] a;
reg [7:0] ld;
reg [7:0] ld2;
reg [7:0] counter [0:50];
reg b = 1'b1;
reg [15:0] x;
reg [5:0] y;

always @(posedge clk or negedge reset) begin
	if (clk | !reset) begin
	if (b) begin
		counter[0] <= 8'b00000000;
		counter[1] <= 8'b00000000;
		counter[2] <= 8'b00000000;
		counter[3] <= 8'b00000000;
		counter[4] <= 8'b00000000;
		counter[5] <= 8'b00000000;
		counter[6] <= 8'b00000000;
		counter[7] <= 8'b00000000;
		counter[8] <= 8'b00000000;
		counter[9] <= 8'b00000000;
		counter[10] <= 8'b00000000;
		counter[11] <= 8'b00000000;
		counter[12] <= 8'b00000000;
		counter[13] <= 8'b00000000;
		counter[14] <= 8'b00000000;
		counter[15] <= 8'b00000000;
		counter[16] <= 8'b00000000;
		counter[17] <= 8'b00000000;
		counter[18] <= 8'b00000000;
		counter[19] <= 8'b00000000;
		counter[20] <= 8'b00000000;
		counter[21] <= 8'b00000000;
		counter[22] <= 8'b00000000;
		counter[23] <= 8'b00000000;
		counter[24] <= 8'b00000000;
		counter[25] <= 8'b00000000;
		counter[26] <= 8'b00000000;
		counter[27] <= 8'b00000000;
		counter[28] <= 8'b00000000;
		counter[29] <= 8'b00000000;
		counter[30] <= 8'b00000000;
		counter[31] <= 8'b00000000;
		counter[32] <= 8'b00000000;
		counter[33] <= 8'b00000000;
		counter[34] <= 8'b00000000;
		counter[35] <= 8'b00000000;
		counter[36] <= 8'b00000000;
		counter[37] <= 8'b00000000;
		counter[38] <= 8'b00000000;
		counter[39] <= 8'b00000000;
		counter[40] <= 8'b00000000;
		counter[41] <= 8'b00000000;
		counter[42] <= 8'b00000000;
		counter[43] <= 8'b00000000;
		counter[44] <= 8'b00000000;
		counter[45] <= 8'b00000000;
		counter[46] <= 8'b00000000;
		counter[47] <= 8'b00000000;
		counter[48] <= 8'b00000000;
		counter[49] <= 8'b00000000;
		counter[50] <= 8'b00000000;
		a <= 10'b0000000000;
		b <= 1'b0;
		x = 16'b0000000000000000;
		y = 6'b000000;
		ld = 8'b00000000;
		ld2 = 8'b00000000; 
	end
	x = x + 16'b0000000000000001;
	case(x)
		16'b0111111111111111: ld2 <= 8'b00000000;
		16'b1111111111111111: begin x = 16'b0000000000000000 ; y = y + 6'b000001 ; ld2 <= counter[y];
			if (y==6'b111111) begin
				y = 6'b000000; end
			end
		default: ; // Default case
	endcase
	if ( signal & a==10'b0000000000) begin
		a <= 10'b0000000001;
	end
	else if ( signal & a!=10'b0000000000) begin
		counter[0] <= counter[0] + 8'b00000001;
		case(a)
			10'b0000000001: counter[1] <= counter[1] + 1;
			10'b0000000010: counter[1] <= counter[1] + 1;
			10'b0000000011: counter[1] <= counter[1] + 1;
			10'b0000000100: counter[1] <= counter[1] + 1;
			10'b0000000101: counter[1] <= counter[1] + 1;
			10'b0000000110: counter[1] <= counter[1] + 1;
			10'b0000000111: counter[1] <= counter[1] + 1;
			10'b0000001000: counter[1] <= counter[1] + 1;
			10'b0000001001: counter[1] <= counter[1] + 1;
			10'b0000001010: counter[1] <= counter[1] + 1;
			10'b0000001011: counter[1] <= counter[1] + 1;
			10'b0000001100: counter[1] <= counter[1] + 1;
			10'b0000001101: counter[1] <= counter[1] + 1;
			10'b0000001110: counter[1] <= counter[1] + 1;
			10'b0000001111: counter[1] <= counter[1] + 1;
			10'b0000010000: counter[1] <= counter[1] + 1;
			10'b0000010001: counter[1] <= counter[1] + 1;
			10'b0000010010: counter[1] <= counter[1] + 1;
			10'b0000010011: counter[1] <= counter[1] + 1;
			10'b0000010100: counter[1] <= counter[1] + 1;
			10'b0000010101: counter[2] <= counter[2] + 1;
			10'b0000010110: counter[2] <= counter[2] + 1;
			10'b0000010111: counter[2] <= counter[2] + 1;
			10'b0000011000: counter[2] <= counter[2] + 1;
			10'b0000011001: counter[2] <= counter[2] + 1;
			10'b0000011010: counter[2] <= counter[2] + 1;
			10'b0000011011: counter[2] <= counter[2] + 1;
			10'b0000011100: counter[2] <= counter[2] + 1;
			10'b0000011101: counter[2] <= counter[2] + 1;
			10'b0000011110: counter[2] <= counter[2] + 1;
			10'b0000011111: counter[2] <= counter[2] + 1;
			10'b0000100000: counter[2] <= counter[2] + 1;
			10'b0000100001: counter[2] <= counter[2] + 1;
			10'b0000100010: counter[2] <= counter[2] + 1;
			10'b0000100011: counter[2] <= counter[2] + 1;
			10'b0000100100: counter[2] <= counter[2] + 1;
			10'b0000100101: counter[2] <= counter[2] + 1;
			10'b0000100110: counter[2] <= counter[2] + 1;
			10'b0000100111: counter[2] <= counter[2] + 1;
			10'b0000101000: counter[2] <= counter[2] + 1;
			10'b0000101001: counter[3] <= counter[3] + 1;
			10'b0000101010: counter[3] <= counter[3] + 1;
			10'b0000101011: counter[3] <= counter[3] + 1;
			10'b0000101100: counter[3] <= counter[3] + 1;
			10'b0000101101: counter[3] <= counter[3] + 1;
			10'b0000101110: counter[3] <= counter[3] + 1;
			10'b0000101111: counter[3] <= counter[3] + 1;
			10'b0000110000: counter[3] <= counter[3] + 1;
			10'b0000110001: counter[3] <= counter[3] + 1;
			10'b0000110010: counter[3] <= counter[3] + 1;
			10'b0000110011: counter[3] <= counter[3] + 1;
			10'b0000110100: counter[3] <= counter[3] + 1;
			10'b0000110101: counter[3] <= counter[3] + 1;
			10'b0000110110: counter[3] <= counter[3] + 1;
			10'b0000110111: counter[3] <= counter[3] + 1;
			10'b0000111000: counter[3] <= counter[3] + 1;
			10'b0000111001: counter[3] <= counter[3] + 1;
			10'b0000111010: counter[3] <= counter[3] + 1;
			10'b0000111011: counter[3] <= counter[3] + 1;
			10'b0000111100: counter[3] <= counter[3] + 1;
			10'b0000111101: counter[4] <= counter[4] + 1;
			10'b0000111110: counter[4] <= counter[4] + 1;
			10'b0000111111: counter[4] <= counter[4] + 1;
			10'b0001000000: counter[4] <= counter[4] + 1;
			10'b0001000001: counter[4] <= counter[4] + 1;
			10'b0001000010: counter[4] <= counter[4] + 1;
			10'b0001000011: counter[4] <= counter[4] + 1;
			10'b0001000100: counter[4] <= counter[4] + 1;
			10'b0001000101: counter[4] <= counter[4] + 1;
			10'b0001000110: counter[4] <= counter[4] + 1;
			10'b0001000111: counter[4] <= counter[4] + 1;
			10'b0001001000: counter[4] <= counter[4] + 1;
			10'b0001001001: counter[4] <= counter[4] + 1;
			10'b0001001010: counter[4] <= counter[4] + 1;
			10'b0001001011: counter[4] <= counter[4] + 1;
			10'b0001001100: counter[4] <= counter[4] + 1;
			10'b0001001101: counter[4] <= counter[4] + 1;
			10'b0001001110: counter[4] <= counter[4] + 1;
			10'b0001001111: counter[4] <= counter[4] + 1;
			10'b0001010000: counter[4] <= counter[4] + 1;
			10'b0001010001: counter[5] <= counter[5] + 1;
			10'b0001010010: counter[5] <= counter[5] + 1;
			10'b0001010011: counter[5] <= counter[5] + 1;
			10'b0001010100: counter[5] <= counter[5] + 1;
			10'b0001010101: counter[5] <= counter[5] + 1;
			10'b0001010110: counter[5] <= counter[5] + 1;
			10'b0001010111: counter[5] <= counter[5] + 1;
			10'b0001011000: counter[5] <= counter[5] + 1;
			10'b0001011001: counter[5] <= counter[5] + 1;
			10'b0001011010: counter[5] <= counter[5] + 1;
			10'b0001011011: counter[5] <= counter[5] + 1;
			10'b0001011100: counter[5] <= counter[5] + 1;
			10'b0001011101: counter[5] <= counter[5] + 1;
			10'b0001011110: counter[5] <= counter[5] + 1;
			10'b0001011111: counter[5] <= counter[5] + 1;
			10'b0001100000: counter[5] <= counter[5] + 1;
			10'b0001100001: counter[5] <= counter[5] + 1;
			10'b0001100010: counter[5] <= counter[5] + 1;
			10'b0001100011: counter[5] <= counter[5] + 1;
			10'b0001100100: counter[5] <= counter[5] + 1;
			10'b0001100101: counter[6] <= counter[6] + 1;
			10'b0001100110: counter[6] <= counter[6] + 1;
			10'b0001100111: counter[6] <= counter[6] + 1;
			10'b0001101000: counter[6] <= counter[6] + 1;
			10'b0001101001: counter[6] <= counter[6] + 1;
			10'b0001101010: counter[6] <= counter[6] + 1;
			10'b0001101011: counter[6] <= counter[6] + 1;
			10'b0001101100: counter[6] <= counter[6] + 1;
			10'b0001101101: counter[6] <= counter[6] + 1;
			10'b0001101110: counter[6] <= counter[6] + 1;
			10'b0001101111: counter[6] <= counter[6] + 1;
			10'b0001110000: counter[6] <= counter[6] + 1;
			10'b0001110001: counter[6] <= counter[6] + 1;
			10'b0001110010: counter[6] <= counter[6] + 1;
			10'b0001110011: counter[6] <= counter[6] + 1;
			10'b0001110100: counter[6] <= counter[6] + 1;
			10'b0001110101: counter[6] <= counter[6] + 1;
			10'b0001110110: counter[6] <= counter[6] + 1;
			10'b0001110111: counter[6] <= counter[6] + 1;
			10'b0001111000: counter[6] <= counter[6] + 1;
			10'b0001111001: counter[7] <= counter[7] + 1;
			10'b0001111010: counter[7] <= counter[7] + 1;
			10'b0001111011: counter[7] <= counter[7] + 1;
			10'b0001111100: counter[7] <= counter[7] + 1;
			10'b0001111101: counter[7] <= counter[7] + 1;
			10'b0001111110: counter[7] <= counter[7] + 1;
			10'b0001111111: counter[7] <= counter[7] + 1;
			10'b0010000000: counter[7] <= counter[7] + 1;
			10'b0010000001: counter[7] <= counter[7] + 1;
			10'b0010000010: counter[7] <= counter[7] + 1;
			10'b0010000011: counter[7] <= counter[7] + 1;
			10'b0010000100: counter[7] <= counter[7] + 1;
			10'b0010000101: counter[7] <= counter[7] + 1;
			10'b0010000110: counter[7] <= counter[7] + 1;
			10'b0010000111: counter[7] <= counter[7] + 1;
			10'b0010001000: counter[7] <= counter[7] + 1;
			10'b0010001001: counter[7] <= counter[7] + 1;
			10'b0010001010: counter[7] <= counter[7] + 1;
			10'b0010001011: counter[7] <= counter[7] + 1;
			10'b0010001100: counter[7] <= counter[7] + 1;
			10'b0010001101: counter[8] <= counter[8] + 1;
			10'b0010001110: counter[8] <= counter[8] + 1;
			10'b0010001111: counter[8] <= counter[8] + 1;
			10'b0010010000: counter[8] <= counter[8] + 1;
			10'b0010010001: counter[8] <= counter[8] + 1;
			10'b0010010010: counter[8] <= counter[8] + 1;
			10'b0010010011: counter[8] <= counter[8] + 1;
			10'b0010010100: counter[8] <= counter[8] + 1;
			10'b0010010101: counter[8] <= counter[8] + 1;
			10'b0010010110: counter[8] <= counter[8] + 1;
			10'b0010010111: counter[8] <= counter[8] + 1;
			10'b0010011000: counter[8] <= counter[8] + 1;
			10'b0010011001: counter[8] <= counter[8] + 1;
			10'b0010011010: counter[8] <= counter[8] + 1;
			10'b0010011011: counter[8] <= counter[8] + 1;
			10'b0010011100: counter[8] <= counter[8] + 1;
			10'b0010011101: counter[8] <= counter[8] + 1;
			10'b0010011110: counter[8] <= counter[8] + 1;
			10'b0010011111: counter[8] <= counter[8] + 1;
			10'b0010100000: counter[8] <= counter[8] + 1;
			10'b0010100001: counter[9] <= counter[9] + 1;
			10'b0010100010: counter[9] <= counter[9] + 1;
			10'b0010100011: counter[9] <= counter[9] + 1;
			10'b0010100100: counter[9] <= counter[9] + 1;
			10'b0010100101: counter[9] <= counter[9] + 1;
			10'b0010100110: counter[9] <= counter[9] + 1;
			10'b0010100111: counter[9] <= counter[9] + 1;
			10'b0010101000: counter[9] <= counter[9] + 1;
			10'b0010101001: counter[9] <= counter[9] + 1;
			10'b0010101010: counter[9] <= counter[9] + 1;
			10'b0010101011: counter[9] <= counter[9] + 1;
			10'b0010101100: counter[9] <= counter[9] + 1;
			10'b0010101101: counter[9] <= counter[9] + 1;
			10'b0010101110: counter[9] <= counter[9] + 1;
			10'b0010101111: counter[9] <= counter[9] + 1;
			10'b0010110000: counter[9] <= counter[9] + 1;
			10'b0010110001: counter[9] <= counter[9] + 1;
			10'b0010110010: counter[9] <= counter[9] + 1;
			10'b0010110011: counter[9] <= counter[9] + 1;
			10'b0010110100: counter[9] <= counter[9] + 1;
			10'b0010110101: counter[10] <= counter[10] + 1;
			10'b0010110110: counter[10] <= counter[10] + 1;
			10'b0010110111: counter[10] <= counter[10] + 1;
			10'b0010111000: counter[10] <= counter[10] + 1;
			10'b0010111001: counter[10] <= counter[10] + 1;
			10'b0010111010: counter[10] <= counter[10] + 1;
			10'b0010111011: counter[10] <= counter[10] + 1;
			10'b0010111100: counter[10] <= counter[10] + 1;
			10'b0010111101: counter[10] <= counter[10] + 1;
			10'b0010111110: counter[10] <= counter[10] + 1;
			10'b0010111111: counter[10] <= counter[10] + 1;
			10'b0011000000: counter[10] <= counter[10] + 1;
			10'b0011000001: counter[10] <= counter[10] + 1;
			10'b0011000010: counter[10] <= counter[10] + 1;
			10'b0011000011: counter[10] <= counter[10] + 1;
			10'b0011000100: counter[10] <= counter[10] + 1;
			10'b0011000101: counter[10] <= counter[10] + 1;
			10'b0011000110: counter[10] <= counter[10] + 1;
			10'b0011000111: counter[10] <= counter[10] + 1;
			10'b0011001000: counter[10] <= counter[10] + 1;
			10'b0011001001: counter[11] <= counter[11] + 1;
			10'b0011001010: counter[11] <= counter[11] + 1;
			10'b0011001011: counter[11] <= counter[11] + 1;
			10'b0011001100: counter[11] <= counter[11] + 1;
			10'b0011001101: counter[11] <= counter[11] + 1;
			10'b0011001110: counter[11] <= counter[11] + 1;
			10'b0011001111: counter[11] <= counter[11] + 1;
			10'b0011010000: counter[11] <= counter[11] + 1;
			10'b0011010001: counter[11] <= counter[11] + 1;
			10'b0011010010: counter[11] <= counter[11] + 1;
			10'b0011010011: counter[11] <= counter[11] + 1;
			10'b0011010100: counter[11] <= counter[11] + 1;
			10'b0011010101: counter[11] <= counter[11] + 1;
			10'b0011010110: counter[11] <= counter[11] + 1;
			10'b0011010111: counter[11] <= counter[11] + 1;
			10'b0011011000: counter[11] <= counter[11] + 1;
			10'b0011011001: counter[11] <= counter[11] + 1;
			10'b0011011010: counter[11] <= counter[11] + 1;
			10'b0011011011: counter[11] <= counter[11] + 1;
			10'b0011011100: counter[11] <= counter[11] + 1;
			10'b0011011101: counter[12] <= counter[12] + 1;
			10'b0011011110: counter[12] <= counter[12] + 1;
			10'b0011011111: counter[12] <= counter[12] + 1;
			10'b0011100000: counter[12] <= counter[12] + 1;
			10'b0011100001: counter[12] <= counter[12] + 1;
			10'b0011100010: counter[12] <= counter[12] + 1;
			10'b0011100011: counter[12] <= counter[12] + 1;
			10'b0011100100: counter[12] <= counter[12] + 1;
			10'b0011100101: counter[12] <= counter[12] + 1;
			10'b0011100110: counter[12] <= counter[12] + 1;
			10'b0011100111: counter[12] <= counter[12] + 1;
			10'b0011101000: counter[12] <= counter[12] + 1;
			10'b0011101001: counter[12] <= counter[12] + 1;
			10'b0011101010: counter[12] <= counter[12] + 1;
			10'b0011101011: counter[12] <= counter[12] + 1;
			10'b0011101100: counter[12] <= counter[12] + 1;
			10'b0011101101: counter[12] <= counter[12] + 1;
			10'b0011101110: counter[12] <= counter[12] + 1;
			10'b0011101111: counter[12] <= counter[12] + 1;
			10'b0011110000: counter[12] <= counter[12] + 1;
			10'b0011110001: counter[13] <= counter[13] + 1;
			10'b0011110010: counter[13] <= counter[13] + 1;
			10'b0011110011: counter[13] <= counter[13] + 1;
			10'b0011110100: counter[13] <= counter[13] + 1;
			10'b0011110101: counter[13] <= counter[13] + 1;
			10'b0011110110: counter[13] <= counter[13] + 1;
			10'b0011110111: counter[13] <= counter[13] + 1;
			10'b0011111000: counter[13] <= counter[13] + 1;
			10'b0011111001: counter[13] <= counter[13] + 1;
			10'b0011111010: counter[13] <= counter[13] + 1;
			10'b0011111011: counter[13] <= counter[13] + 1;
			10'b0011111100: counter[13] <= counter[13] + 1;
			10'b0011111101: counter[13] <= counter[13] + 1;
			10'b0011111110: counter[13] <= counter[13] + 1;
			10'b0011111111: counter[13] <= counter[13] + 1;
			10'b0100000000: counter[13] <= counter[13] + 1;
			10'b0100000001: counter[13] <= counter[13] + 1;
			10'b0100000010: counter[13] <= counter[13] + 1;
			10'b0100000011: counter[13] <= counter[13] + 1;
			10'b0100000100: counter[13] <= counter[13] + 1;
			10'b0100000101: counter[14] <= counter[14] + 1;
			10'b0100000110: counter[14] <= counter[14] + 1;
			10'b0100000111: counter[14] <= counter[14] + 1;
			10'b0100001000: counter[14] <= counter[14] + 1;
			10'b0100001001: counter[14] <= counter[14] + 1;
			10'b0100001010: counter[14] <= counter[14] + 1;
			10'b0100001011: counter[14] <= counter[14] + 1;
			10'b0100001100: counter[14] <= counter[14] + 1;
			10'b0100001101: counter[14] <= counter[14] + 1;
			10'b0100001110: counter[14] <= counter[14] + 1;
			10'b0100001111: counter[14] <= counter[14] + 1;
			10'b0100010000: counter[14] <= counter[14] + 1;
			10'b0100010001: counter[14] <= counter[14] + 1;
			10'b0100010010: counter[14] <= counter[14] + 1;
			10'b0100010011: counter[14] <= counter[14] + 1;
			10'b0100010100: counter[14] <= counter[14] + 1;
			10'b0100010101: counter[14] <= counter[14] + 1;
			10'b0100010110: counter[14] <= counter[14] + 1;
			10'b0100010111: counter[14] <= counter[14] + 1;
			10'b0100011000: counter[14] <= counter[14] + 1;
			10'b0100011001: counter[15] <= counter[15] + 1;
			10'b0100011010: counter[15] <= counter[15] + 1;
			10'b0100011011: counter[15] <= counter[15] + 1;
			10'b0100011100: counter[15] <= counter[15] + 1;
			10'b0100011101: counter[15] <= counter[15] + 1;
			10'b0100011110: counter[15] <= counter[15] + 1;
			10'b0100011111: counter[15] <= counter[15] + 1;
			10'b0100100000: counter[15] <= counter[15] + 1;
			10'b0100100001: counter[15] <= counter[15] + 1;
			10'b0100100010: counter[15] <= counter[15] + 1;
			10'b0100100011: counter[15] <= counter[15] + 1;
			10'b0100100100: counter[15] <= counter[15] + 1;
			10'b0100100101: counter[15] <= counter[15] + 1;
			10'b0100100110: counter[15] <= counter[15] + 1;
			10'b0100100111: counter[15] <= counter[15] + 1;
			10'b0100101000: counter[15] <= counter[15] + 1;
			10'b0100101001: counter[15] <= counter[15] + 1;
			10'b0100101010: counter[15] <= counter[15] + 1;
			10'b0100101011: counter[15] <= counter[15] + 1;
			10'b0100101100: counter[15] <= counter[15] + 1;
			10'b0100101101: counter[16] <= counter[16] + 1;
			10'b0100101110: counter[16] <= counter[16] + 1;
			10'b0100101111: counter[16] <= counter[16] + 1;
			10'b0100110000: counter[16] <= counter[16] + 1;
			10'b0100110001: counter[16] <= counter[16] + 1;
			10'b0100110010: counter[16] <= counter[16] + 1;
			10'b0100110011: counter[16] <= counter[16] + 1;
			10'b0100110100: counter[16] <= counter[16] + 1;
			10'b0100110101: counter[16] <= counter[16] + 1;
			10'b0100110110: counter[16] <= counter[16] + 1;
			10'b0100110111: counter[16] <= counter[16] + 1;
			10'b0100111000: counter[16] <= counter[16] + 1;
			10'b0100111001: counter[16] <= counter[16] + 1;
			10'b0100111010: counter[16] <= counter[16] + 1;
			10'b0100111011: counter[16] <= counter[16] + 1;
			10'b0100111100: counter[16] <= counter[16] + 1;
			10'b0100111101: counter[16] <= counter[16] + 1;
			10'b0100111110: counter[16] <= counter[16] + 1;
			10'b0100111111: counter[16] <= counter[16] + 1;
			10'b0101000000: counter[16] <= counter[16] + 1;
			10'b0101000001: counter[17] <= counter[17] + 1;
			10'b0101000010: counter[17] <= counter[17] + 1;
			10'b0101000011: counter[17] <= counter[17] + 1;
			10'b0101000100: counter[17] <= counter[17] + 1;
			10'b0101000101: counter[17] <= counter[17] + 1;
			10'b0101000110: counter[17] <= counter[17] + 1;
			10'b0101000111: counter[17] <= counter[17] + 1;
			10'b0101001000: counter[17] <= counter[17] + 1;
			10'b0101001001: counter[17] <= counter[17] + 1;
			10'b0101001010: counter[17] <= counter[17] + 1;
			10'b0101001011: counter[17] <= counter[17] + 1;
			10'b0101001100: counter[17] <= counter[17] + 1;
			10'b0101001101: counter[17] <= counter[17] + 1;
			10'b0101001110: counter[17] <= counter[17] + 1;
			10'b0101001111: counter[17] <= counter[17] + 1;
			10'b0101010000: counter[17] <= counter[17] + 1;
			10'b0101010001: counter[17] <= counter[17] + 1;
			10'b0101010010: counter[17] <= counter[17] + 1;
			10'b0101010011: counter[17] <= counter[17] + 1;
			10'b0101010100: counter[17] <= counter[17] + 1;
			10'b0101010101: counter[18] <= counter[18] + 1;
			10'b0101010110: counter[18] <= counter[18] + 1;
			10'b0101010111: counter[18] <= counter[18] + 1;
			10'b0101011000: counter[18] <= counter[18] + 1;
			10'b0101011001: counter[18] <= counter[18] + 1;
			10'b0101011010: counter[18] <= counter[18] + 1;
			10'b0101011011: counter[18] <= counter[18] + 1;
			10'b0101011100: counter[18] <= counter[18] + 1;
			10'b0101011101: counter[18] <= counter[18] + 1;
			10'b0101011110: counter[18] <= counter[18] + 1;
			10'b0101011111: counter[18] <= counter[18] + 1;
			10'b0101100000: counter[18] <= counter[18] + 1;
			10'b0101100001: counter[18] <= counter[18] + 1;
			10'b0101100010: counter[18] <= counter[18] + 1;
			10'b0101100011: counter[18] <= counter[18] + 1;
			10'b0101100100: counter[18] <= counter[18] + 1;
			10'b0101100101: counter[18] <= counter[18] + 1;
			10'b0101100110: counter[18] <= counter[18] + 1;
			10'b0101100111: counter[18] <= counter[18] + 1;
			10'b0101101000: counter[18] <= counter[18] + 1;
			10'b0101101001: counter[19] <= counter[19] + 1;
			10'b0101101010: counter[19] <= counter[19] + 1;
			10'b0101101011: counter[19] <= counter[19] + 1;
			10'b0101101100: counter[19] <= counter[19] + 1;
			10'b0101101101: counter[19] <= counter[19] + 1;
			10'b0101101110: counter[19] <= counter[19] + 1;
			10'b0101101111: counter[19] <= counter[19] + 1;
			10'b0101110000: counter[19] <= counter[19] + 1;
			10'b0101110001: counter[19] <= counter[19] + 1;
			10'b0101110010: counter[19] <= counter[19] + 1;
			10'b0101110011: counter[19] <= counter[19] + 1;
			10'b0101110100: counter[19] <= counter[19] + 1;
			10'b0101110101: counter[19] <= counter[19] + 1;
			10'b0101110110: counter[19] <= counter[19] + 1;
			10'b0101110111: counter[19] <= counter[19] + 1;
			10'b0101111000: counter[19] <= counter[19] + 1;
			10'b0101111001: counter[19] <= counter[19] + 1;
			10'b0101111010: counter[19] <= counter[19] + 1;
			10'b0101111011: counter[19] <= counter[19] + 1;
			10'b0101111100: counter[19] <= counter[19] + 1;
			10'b0101111101: counter[20] <= counter[20] + 1;
			10'b0101111110: counter[20] <= counter[20] + 1;
			10'b0101111111: counter[20] <= counter[20] + 1;
			10'b0110000000: counter[20] <= counter[20] + 1;
			10'b0110000001: counter[20] <= counter[20] + 1;
			10'b0110000010: counter[20] <= counter[20] + 1;
			10'b0110000011: counter[20] <= counter[20] + 1;
			10'b0110000100: counter[20] <= counter[20] + 1;
			10'b0110000101: counter[20] <= counter[20] + 1;
			10'b0110000110: counter[20] <= counter[20] + 1;
			10'b0110000111: counter[20] <= counter[20] + 1;
			10'b0110001000: counter[20] <= counter[20] + 1;
			10'b0110001001: counter[20] <= counter[20] + 1;
			10'b0110001010: counter[20] <= counter[20] + 1;
			10'b0110001011: counter[20] <= counter[20] + 1;
			10'b0110001100: counter[20] <= counter[20] + 1;
			10'b0110001101: counter[20] <= counter[20] + 1;
			10'b0110001110: counter[20] <= counter[20] + 1;
			10'b0110001111: counter[20] <= counter[20] + 1;
			10'b0110010000: counter[20] <= counter[20] + 1;
			10'b0110010001: counter[21] <= counter[21] + 1;
			10'b0110010010: counter[21] <= counter[21] + 1;
			10'b0110010011: counter[21] <= counter[21] + 1;
			10'b0110010100: counter[21] <= counter[21] + 1;
			10'b0110010101: counter[21] <= counter[21] + 1;
			10'b0110010110: counter[21] <= counter[21] + 1;
			10'b0110010111: counter[21] <= counter[21] + 1;
			10'b0110011000: counter[21] <= counter[21] + 1;
			10'b0110011001: counter[21] <= counter[21] + 1;
			10'b0110011010: counter[21] <= counter[21] + 1;
			10'b0110011011: counter[21] <= counter[21] + 1;
			10'b0110011100: counter[21] <= counter[21] + 1;
			10'b0110011101: counter[21] <= counter[21] + 1;
			10'b0110011110: counter[21] <= counter[21] + 1;
			10'b0110011111: counter[21] <= counter[21] + 1;
			10'b0110100000: counter[21] <= counter[21] + 1;
			10'b0110100001: counter[21] <= counter[21] + 1;
			10'b0110100010: counter[21] <= counter[21] + 1;
			10'b0110100011: counter[21] <= counter[21] + 1;
			10'b0110100100: counter[21] <= counter[21] + 1;
			10'b0110100101: counter[22] <= counter[22] + 1;
			10'b0110100110: counter[22] <= counter[22] + 1;
			10'b0110100111: counter[22] <= counter[22] + 1;
			10'b0110101000: counter[22] <= counter[22] + 1;
			10'b0110101001: counter[22] <= counter[22] + 1;
			10'b0110101010: counter[22] <= counter[22] + 1;
			10'b0110101011: counter[22] <= counter[22] + 1;
			10'b0110101100: counter[22] <= counter[22] + 1;
			10'b0110101101: counter[22] <= counter[22] + 1;
			10'b0110101110: counter[22] <= counter[22] + 1;
			10'b0110101111: counter[22] <= counter[22] + 1;
			10'b0110110000: counter[22] <= counter[22] + 1;
			10'b0110110001: counter[22] <= counter[22] + 1;
			10'b0110110010: counter[22] <= counter[22] + 1;
			10'b0110110011: counter[22] <= counter[22] + 1;
			10'b0110110100: counter[22] <= counter[22] + 1;
			10'b0110110101: counter[22] <= counter[22] + 1;
			10'b0110110110: counter[22] <= counter[22] + 1;
			10'b0110110111: counter[22] <= counter[22] + 1;
			10'b0110111000: counter[22] <= counter[22] + 1;
			10'b0110111001: counter[23] <= counter[23] + 1;
			10'b0110111010: counter[23] <= counter[23] + 1;
			10'b0110111011: counter[23] <= counter[23] + 1;
			10'b0110111100: counter[23] <= counter[23] + 1;
			10'b0110111101: counter[23] <= counter[23] + 1;
			10'b0110111110: counter[23] <= counter[23] + 1;
			10'b0110111111: counter[23] <= counter[23] + 1;
			10'b0111000000: counter[23] <= counter[23] + 1;
			10'b0111000001: counter[23] <= counter[23] + 1;
			10'b0111000010: counter[23] <= counter[23] + 1;
			10'b0111000011: counter[23] <= counter[23] + 1;
			10'b0111000100: counter[23] <= counter[23] + 1;
			10'b0111000101: counter[23] <= counter[23] + 1;
			10'b0111000110: counter[23] <= counter[23] + 1;
			10'b0111000111: counter[23] <= counter[23] + 1;
			10'b0111001000: counter[23] <= counter[23] + 1;
			10'b0111001001: counter[23] <= counter[23] + 1;
			10'b0111001010: counter[23] <= counter[23] + 1;
			10'b0111001011: counter[23] <= counter[23] + 1;
			10'b0111001100: counter[23] <= counter[23] + 1;
			10'b0111001101: counter[24] <= counter[24] + 1;
			10'b0111001110: counter[24] <= counter[24] + 1;
			10'b0111001111: counter[24] <= counter[24] + 1;
			10'b0111010000: counter[24] <= counter[24] + 1;
			10'b0111010001: counter[24] <= counter[24] + 1;
			10'b0111010010: counter[24] <= counter[24] + 1;
			10'b0111010011: counter[24] <= counter[24] + 1;
			10'b0111010100: counter[24] <= counter[24] + 1;
			10'b0111010101: counter[24] <= counter[24] + 1;
			10'b0111010110: counter[24] <= counter[24] + 1;
			10'b0111010111: counter[24] <= counter[24] + 1;
			10'b0111011000: counter[24] <= counter[24] + 1;
			10'b0111011001: counter[24] <= counter[24] + 1;
			10'b0111011010: counter[24] <= counter[24] + 1;
			10'b0111011011: counter[24] <= counter[24] + 1;
			10'b0111011100: counter[24] <= counter[24] + 1;
			10'b0111011101: counter[24] <= counter[24] + 1;
			10'b0111011110: counter[24] <= counter[24] + 1;
			10'b0111011111: counter[24] <= counter[24] + 1;
			10'b0111100000: counter[24] <= counter[24] + 1;
			10'b0111100001: counter[25] <= counter[25] + 1;
			10'b0111100010: counter[25] <= counter[25] + 1;
			10'b0111100011: counter[25] <= counter[25] + 1;
			10'b0111100100: counter[25] <= counter[25] + 1;
			10'b0111100101: counter[25] <= counter[25] + 1;
			10'b0111100110: counter[25] <= counter[25] + 1;
			10'b0111100111: counter[25] <= counter[25] + 1;
			10'b0111101000: counter[25] <= counter[25] + 1;
			10'b0111101001: counter[25] <= counter[25] + 1;
			10'b0111101010: counter[25] <= counter[25] + 1;
			10'b0111101011: counter[25] <= counter[25] + 1;
			10'b0111101100: counter[25] <= counter[25] + 1;
			10'b0111101101: counter[25] <= counter[25] + 1;
			10'b0111101110: counter[25] <= counter[25] + 1;
			10'b0111101111: counter[25] <= counter[25] + 1;
			10'b0111110000: counter[25] <= counter[25] + 1;
			10'b0111110001: counter[25] <= counter[25] + 1;
			10'b0111110010: counter[25] <= counter[25] + 1;
			10'b0111110011: counter[25] <= counter[25] + 1;
			10'b0111110100: counter[25] <= counter[25] + 1;
			10'b0111110101: counter[26] <= counter[26] + 1;
			10'b0111110110: counter[26] <= counter[26] + 1;
			10'b0111110111: counter[26] <= counter[26] + 1;
			10'b0111111000: counter[26] <= counter[26] + 1;
			10'b0111111001: counter[26] <= counter[26] + 1;
			10'b0111111010: counter[26] <= counter[26] + 1;
			10'b0111111011: counter[26] <= counter[26] + 1;
			10'b0111111100: counter[26] <= counter[26] + 1;
			10'b0111111101: counter[26] <= counter[26] + 1;
			10'b0111111110: counter[26] <= counter[26] + 1;
			10'b0111111111: counter[26] <= counter[26] + 1;
			10'b1000000000: counter[26] <= counter[26] + 1;
			10'b1000000001: counter[26] <= counter[26] + 1;
			10'b1000000010: counter[26] <= counter[26] + 1;
			10'b1000000011: counter[26] <= counter[26] + 1;
			10'b1000000100: counter[26] <= counter[26] + 1;
			10'b1000000101: counter[26] <= counter[26] + 1;
			10'b1000000110: counter[26] <= counter[26] + 1;
			10'b1000000111: counter[26] <= counter[26] + 1;
			10'b1000001000: counter[26] <= counter[26] + 1;
			10'b1000001001: counter[27] <= counter[27] + 1;
			10'b1000001010: counter[27] <= counter[27] + 1;
			10'b1000001011: counter[27] <= counter[27] + 1;
			10'b1000001100: counter[27] <= counter[27] + 1;
			10'b1000001101: counter[27] <= counter[27] + 1;
			10'b1000001110: counter[27] <= counter[27] + 1;
			10'b1000001111: counter[27] <= counter[27] + 1;
			10'b1000010000: counter[27] <= counter[27] + 1;
			10'b1000010001: counter[27] <= counter[27] + 1;
			10'b1000010010: counter[27] <= counter[27] + 1;
			10'b1000010011: counter[27] <= counter[27] + 1;
			10'b1000010100: counter[27] <= counter[27] + 1;
			10'b1000010101: counter[27] <= counter[27] + 1;
			10'b1000010110: counter[27] <= counter[27] + 1;
			10'b1000010111: counter[27] <= counter[27] + 1;
			10'b1000011000: counter[27] <= counter[27] + 1;
			10'b1000011001: counter[27] <= counter[27] + 1;
			10'b1000011010: counter[27] <= counter[27] + 1;
			10'b1000011011: counter[27] <= counter[27] + 1;
			10'b1000011100: counter[27] <= counter[27] + 1;
			10'b1000011101: counter[28] <= counter[28] + 1;
			10'b1000011110: counter[28] <= counter[28] + 1;
			10'b1000011111: counter[28] <= counter[28] + 1;
			10'b1000100000: counter[28] <= counter[28] + 1;
			10'b1000100001: counter[28] <= counter[28] + 1;
			10'b1000100010: counter[28] <= counter[28] + 1;
			10'b1000100011: counter[28] <= counter[28] + 1;
			10'b1000100100: counter[28] <= counter[28] + 1;
			10'b1000100101: counter[28] <= counter[28] + 1;
			10'b1000100110: counter[28] <= counter[28] + 1;
			10'b1000100111: counter[28] <= counter[28] + 1;
			10'b1000101000: counter[28] <= counter[28] + 1;
			10'b1000101001: counter[28] <= counter[28] + 1;
			10'b1000101010: counter[28] <= counter[28] + 1;
			10'b1000101011: counter[28] <= counter[28] + 1;
			10'b1000101100: counter[28] <= counter[28] + 1;
			10'b1000101101: counter[28] <= counter[28] + 1;
			10'b1000101110: counter[28] <= counter[28] + 1;
			10'b1000101111: counter[28] <= counter[28] + 1;
			10'b1000110000: counter[28] <= counter[28] + 1;
			10'b1000110001: counter[29] <= counter[29] + 1;
			10'b1000110010: counter[29] <= counter[29] + 1;
			10'b1000110011: counter[29] <= counter[29] + 1;
			10'b1000110100: counter[29] <= counter[29] + 1;
			10'b1000110101: counter[29] <= counter[29] + 1;
			10'b1000110110: counter[29] <= counter[29] + 1;
			10'b1000110111: counter[29] <= counter[29] + 1;
			10'b1000111000: counter[29] <= counter[29] + 1;
			10'b1000111001: counter[29] <= counter[29] + 1;
			10'b1000111010: counter[29] <= counter[29] + 1;
			10'b1000111011: counter[29] <= counter[29] + 1;
			10'b1000111100: counter[29] <= counter[29] + 1;
			10'b1000111101: counter[29] <= counter[29] + 1;
			10'b1000111110: counter[29] <= counter[29] + 1;
			10'b1000111111: counter[29] <= counter[29] + 1;
			10'b1001000000: counter[29] <= counter[29] + 1;
			10'b1001000001: counter[29] <= counter[29] + 1;
			10'b1001000010: counter[29] <= counter[29] + 1;
			10'b1001000011: counter[29] <= counter[29] + 1;
			10'b1001000100: counter[29] <= counter[29] + 1;
			10'b1001000101: counter[30] <= counter[30] + 1;
			10'b1001000110: counter[30] <= counter[30] + 1;
			10'b1001000111: counter[30] <= counter[30] + 1;
			10'b1001001000: counter[30] <= counter[30] + 1;
			10'b1001001001: counter[30] <= counter[30] + 1;
			10'b1001001010: counter[30] <= counter[30] + 1;
			10'b1001001011: counter[30] <= counter[30] + 1;
			10'b1001001100: counter[30] <= counter[30] + 1;
			10'b1001001101: counter[30] <= counter[30] + 1;
			10'b1001001110: counter[30] <= counter[30] + 1;
			10'b1001001111: counter[30] <= counter[30] + 1;
			10'b1001010000: counter[30] <= counter[30] + 1;
			10'b1001010001: counter[30] <= counter[30] + 1;
			10'b1001010010: counter[30] <= counter[30] + 1;
			10'b1001010011: counter[30] <= counter[30] + 1;
			10'b1001010100: counter[30] <= counter[30] + 1;
			10'b1001010101: counter[30] <= counter[30] + 1;
			10'b1001010110: counter[30] <= counter[30] + 1;
			10'b1001010111: counter[30] <= counter[30] + 1;
			10'b1001011000: counter[30] <= counter[30] + 1;
			10'b1001011001: counter[31] <= counter[31] + 1;
			10'b1001011010: counter[31] <= counter[31] + 1;
			10'b1001011011: counter[31] <= counter[31] + 1;
			10'b1001011100: counter[31] <= counter[31] + 1;
			10'b1001011101: counter[31] <= counter[31] + 1;
			10'b1001011110: counter[31] <= counter[31] + 1;
			10'b1001011111: counter[31] <= counter[31] + 1;
			10'b1001100000: counter[31] <= counter[31] + 1;
			10'b1001100001: counter[31] <= counter[31] + 1;
			10'b1001100010: counter[31] <= counter[31] + 1;
			10'b1001100011: counter[31] <= counter[31] + 1;
			10'b1001100100: counter[31] <= counter[31] + 1;
			10'b1001100101: counter[31] <= counter[31] + 1;
			10'b1001100110: counter[31] <= counter[31] + 1;
			10'b1001100111: counter[31] <= counter[31] + 1;
			10'b1001101000: counter[31] <= counter[31] + 1;
			10'b1001101001: counter[31] <= counter[31] + 1;
			10'b1001101010: counter[31] <= counter[31] + 1;
			10'b1001101011: counter[31] <= counter[31] + 1;
			10'b1001101100: counter[31] <= counter[31] + 1;
			10'b1001101101: counter[32] <= counter[32] + 1;
			10'b1001101110: counter[32] <= counter[32] + 1;
			10'b1001101111: counter[32] <= counter[32] + 1;
			10'b1001110000: counter[32] <= counter[32] + 1;
			10'b1001110001: counter[32] <= counter[32] + 1;
			10'b1001110010: counter[32] <= counter[32] + 1;
			10'b1001110011: counter[32] <= counter[32] + 1;
			10'b1001110100: counter[32] <= counter[32] + 1;
			10'b1001110101: counter[32] <= counter[32] + 1;
			10'b1001110110: counter[32] <= counter[32] + 1;
			10'b1001110111: counter[32] <= counter[32] + 1;
			10'b1001111000: counter[32] <= counter[32] + 1;
			10'b1001111001: counter[32] <= counter[32] + 1;
			10'b1001111010: counter[32] <= counter[32] + 1;
			10'b1001111011: counter[32] <= counter[32] + 1;
			10'b1001111100: counter[32] <= counter[32] + 1;
			10'b1001111101: counter[32] <= counter[32] + 1;
			10'b1001111110: counter[32] <= counter[32] + 1;
			10'b1001111111: counter[32] <= counter[32] + 1;
			10'b1010000000: counter[32] <= counter[32] + 1;
			10'b1010000001: counter[33] <= counter[33] + 1;
			10'b1010000010: counter[33] <= counter[33] + 1;
			10'b1010000011: counter[33] <= counter[33] + 1;
			10'b1010000100: counter[33] <= counter[33] + 1;
			10'b1010000101: counter[33] <= counter[33] + 1;
			10'b1010000110: counter[33] <= counter[33] + 1;
			10'b1010000111: counter[33] <= counter[33] + 1;
			10'b1010001000: counter[33] <= counter[33] + 1;
			10'b1010001001: counter[33] <= counter[33] + 1;
			10'b1010001010: counter[33] <= counter[33] + 1;
			10'b1010001011: counter[33] <= counter[33] + 1;
			10'b1010001100: counter[33] <= counter[33] + 1;
			10'b1010001101: counter[33] <= counter[33] + 1;
			10'b1010001110: counter[33] <= counter[33] + 1;
			10'b1010001111: counter[33] <= counter[33] + 1;
			10'b1010010000: counter[33] <= counter[33] + 1;
			10'b1010010001: counter[33] <= counter[33] + 1;
			10'b1010010010: counter[33] <= counter[33] + 1;
			10'b1010010011: counter[33] <= counter[33] + 1;
			10'b1010010100: counter[33] <= counter[33] + 1;
			10'b1010010101: counter[34] <= counter[34] + 1;
			10'b1010010110: counter[34] <= counter[34] + 1;
			10'b1010010111: counter[34] <= counter[34] + 1;
			10'b1010011000: counter[34] <= counter[34] + 1;
			10'b1010011001: counter[34] <= counter[34] + 1;
			10'b1010011010: counter[34] <= counter[34] + 1;
			10'b1010011011: counter[34] <= counter[34] + 1;
			10'b1010011100: counter[34] <= counter[34] + 1;
			10'b1010011101: counter[34] <= counter[34] + 1;
			10'b1010011110: counter[34] <= counter[34] + 1;
			10'b1010011111: counter[34] <= counter[34] + 1;
			10'b1010100000: counter[34] <= counter[34] + 1;
			10'b1010100001: counter[34] <= counter[34] + 1;
			10'b1010100010: counter[34] <= counter[34] + 1;
			10'b1010100011: counter[34] <= counter[34] + 1;
			10'b1010100100: counter[34] <= counter[34] + 1;
			10'b1010100101: counter[34] <= counter[34] + 1;
			10'b1010100110: counter[34] <= counter[34] + 1;
			10'b1010100111: counter[34] <= counter[34] + 1;
			10'b1010101000: counter[34] <= counter[34] + 1;
			10'b1010101001: counter[35] <= counter[35] + 1;
			10'b1010101010: counter[35] <= counter[35] + 1;
			10'b1010101011: counter[35] <= counter[35] + 1;
			10'b1010101100: counter[35] <= counter[35] + 1;
			10'b1010101101: counter[35] <= counter[35] + 1;
			10'b1010101110: counter[35] <= counter[35] + 1;
			10'b1010101111: counter[35] <= counter[35] + 1;
			10'b1010110000: counter[35] <= counter[35] + 1;
			10'b1010110001: counter[35] <= counter[35] + 1;
			10'b1010110010: counter[35] <= counter[35] + 1;
			10'b1010110011: counter[35] <= counter[35] + 1;
			10'b1010110100: counter[35] <= counter[35] + 1;
			10'b1010110101: counter[35] <= counter[35] + 1;
			10'b1010110110: counter[35] <= counter[35] + 1;
			10'b1010110111: counter[35] <= counter[35] + 1;
			10'b1010111000: counter[35] <= counter[35] + 1;
			10'b1010111001: counter[35] <= counter[35] + 1;
			10'b1010111010: counter[35] <= counter[35] + 1;
			10'b1010111011: counter[35] <= counter[35] + 1;
			10'b1010111100: counter[35] <= counter[35] + 1;
			10'b1010111101: counter[36] <= counter[36] + 1;
			10'b1010111110: counter[36] <= counter[36] + 1;
			10'b1010111111: counter[36] <= counter[36] + 1;
			10'b1011000000: counter[36] <= counter[36] + 1;
			10'b1011000001: counter[36] <= counter[36] + 1;
			10'b1011000010: counter[36] <= counter[36] + 1;
			10'b1011000011: counter[36] <= counter[36] + 1;
			10'b1011000100: counter[36] <= counter[36] + 1;
			10'b1011000101: counter[36] <= counter[36] + 1;
			10'b1011000110: counter[36] <= counter[36] + 1;
			10'b1011000111: counter[36] <= counter[36] + 1;
			10'b1011001000: counter[36] <= counter[36] + 1;
			10'b1011001001: counter[36] <= counter[36] + 1;
			10'b1011001010: counter[36] <= counter[36] + 1;
			10'b1011001011: counter[36] <= counter[36] + 1;
			10'b1011001100: counter[36] <= counter[36] + 1;
			10'b1011001101: counter[36] <= counter[36] + 1;
			10'b1011001110: counter[36] <= counter[36] + 1;
			10'b1011001111: counter[36] <= counter[36] + 1;
			10'b1011010000: counter[36] <= counter[36] + 1;
			10'b1011010001: counter[37] <= counter[37] + 1;
			10'b1011010010: counter[37] <= counter[37] + 1;
			10'b1011010011: counter[37] <= counter[37] + 1;
			10'b1011010100: counter[37] <= counter[37] + 1;
			10'b1011010101: counter[37] <= counter[37] + 1;
			10'b1011010110: counter[37] <= counter[37] + 1;
			10'b1011010111: counter[37] <= counter[37] + 1;
			10'b1011011000: counter[37] <= counter[37] + 1;
			10'b1011011001: counter[37] <= counter[37] + 1;
			10'b1011011010: counter[37] <= counter[37] + 1;
			10'b1011011011: counter[37] <= counter[37] + 1;
			10'b1011011100: counter[37] <= counter[37] + 1;
			10'b1011011101: counter[37] <= counter[37] + 1;
			10'b1011011110: counter[37] <= counter[37] + 1;
			10'b1011011111: counter[37] <= counter[37] + 1;
			10'b1011100000: counter[37] <= counter[37] + 1;
			10'b1011100001: counter[37] <= counter[37] + 1;
			10'b1011100010: counter[37] <= counter[37] + 1;
			10'b1011100011: counter[37] <= counter[37] + 1;
			10'b1011100100: counter[37] <= counter[37] + 1;
			10'b1011100101: counter[38] <= counter[38] + 1;
			10'b1011100110: counter[38] <= counter[38] + 1;
			10'b1011100111: counter[38] <= counter[38] + 1;
			10'b1011101000: counter[38] <= counter[38] + 1;
			10'b1011101001: counter[38] <= counter[38] + 1;
			10'b1011101010: counter[38] <= counter[38] + 1;
			10'b1011101011: counter[38] <= counter[38] + 1;
			10'b1011101100: counter[38] <= counter[38] + 1;
			10'b1011101101: counter[38] <= counter[38] + 1;
			10'b1011101110: counter[38] <= counter[38] + 1;
			10'b1011101111: counter[38] <= counter[38] + 1;
			10'b1011110000: counter[38] <= counter[38] + 1;
			10'b1011110001: counter[38] <= counter[38] + 1;
			10'b1011110010: counter[38] <= counter[38] + 1;
			10'b1011110011: counter[38] <= counter[38] + 1;
			10'b1011110100: counter[38] <= counter[38] + 1;
			10'b1011110101: counter[38] <= counter[38] + 1;
			10'b1011110110: counter[38] <= counter[38] + 1;
			10'b1011110111: counter[38] <= counter[38] + 1;
			10'b1011111000: counter[38] <= counter[38] + 1;
			10'b1011111001: counter[39] <= counter[39] + 1;
			10'b1011111010: counter[39] <= counter[39] + 1;
			10'b1011111011: counter[39] <= counter[39] + 1;
			10'b1011111100: counter[39] <= counter[39] + 1;
			10'b1011111101: counter[39] <= counter[39] + 1;
			10'b1011111110: counter[39] <= counter[39] + 1;
			10'b1011111111: counter[39] <= counter[39] + 1;
			10'b1100000000: counter[39] <= counter[39] + 1;
			10'b1100000001: counter[39] <= counter[39] + 1;
			10'b1100000010: counter[39] <= counter[39] + 1;
			10'b1100000011: counter[39] <= counter[39] + 1;
			10'b1100000100: counter[39] <= counter[39] + 1;
			10'b1100000101: counter[39] <= counter[39] + 1;
			10'b1100000110: counter[39] <= counter[39] + 1;
			10'b1100000111: counter[39] <= counter[39] + 1;
			10'b1100001000: counter[39] <= counter[39] + 1;
			10'b1100001001: counter[39] <= counter[39] + 1;
			10'b1100001010: counter[39] <= counter[39] + 1;
			10'b1100001011: counter[39] <= counter[39] + 1;
			10'b1100001100: counter[39] <= counter[39] + 1;
			10'b1100001101: counter[40] <= counter[40] + 1;
			10'b1100001110: counter[40] <= counter[40] + 1;
			10'b1100001111: counter[40] <= counter[40] + 1;
			10'b1100010000: counter[40] <= counter[40] + 1;
			10'b1100010001: counter[40] <= counter[40] + 1;
			10'b1100010010: counter[40] <= counter[40] + 1;
			10'b1100010011: counter[40] <= counter[40] + 1;
			10'b1100010100: counter[40] <= counter[40] + 1;
			10'b1100010101: counter[40] <= counter[40] + 1;
			10'b1100010110: counter[40] <= counter[40] + 1;
			10'b1100010111: counter[40] <= counter[40] + 1;
			10'b1100011000: counter[40] <= counter[40] + 1;
			10'b1100011001: counter[40] <= counter[40] + 1;
			10'b1100011010: counter[40] <= counter[40] + 1;
			10'b1100011011: counter[40] <= counter[40] + 1;
			10'b1100011100: counter[40] <= counter[40] + 1;
			10'b1100011101: counter[40] <= counter[40] + 1;
			10'b1100011110: counter[40] <= counter[40] + 1;
			10'b1100011111: counter[40] <= counter[40] + 1;
			10'b1100100000: counter[40] <= counter[40] + 1;
			10'b1100100001: counter[41] <= counter[41] + 1;
			10'b1100100010: counter[41] <= counter[41] + 1;
			10'b1100100011: counter[41] <= counter[41] + 1;
			10'b1100100100: counter[41] <= counter[41] + 1;
			10'b1100100101: counter[41] <= counter[41] + 1;
			10'b1100100110: counter[41] <= counter[41] + 1;
			10'b1100100111: counter[41] <= counter[41] + 1;
			10'b1100101000: counter[41] <= counter[41] + 1;
			10'b1100101001: counter[41] <= counter[41] + 1;
			10'b1100101010: counter[41] <= counter[41] + 1;
			10'b1100101011: counter[41] <= counter[41] + 1;
			10'b1100101100: counter[41] <= counter[41] + 1;
			10'b1100101101: counter[41] <= counter[41] + 1;
			10'b1100101110: counter[41] <= counter[41] + 1;
			10'b1100101111: counter[41] <= counter[41] + 1;
			10'b1100110000: counter[41] <= counter[41] + 1;
			10'b1100110001: counter[41] <= counter[41] + 1;
			10'b1100110010: counter[41] <= counter[41] + 1;
			10'b1100110011: counter[41] <= counter[41] + 1;
			10'b1100110100: counter[41] <= counter[41] + 1;
			10'b1100110101: counter[42] <= counter[42] + 1;
			10'b1100110110: counter[42] <= counter[42] + 1;
			10'b1100110111: counter[42] <= counter[42] + 1;
			10'b1100111000: counter[42] <= counter[42] + 1;
			10'b1100111001: counter[42] <= counter[42] + 1;
			10'b1100111010: counter[42] <= counter[42] + 1;
			10'b1100111011: counter[42] <= counter[42] + 1;
			10'b1100111100: counter[42] <= counter[42] + 1;
			10'b1100111101: counter[42] <= counter[42] + 1;
			10'b1100111110: counter[42] <= counter[42] + 1;
			10'b1100111111: counter[42] <= counter[42] + 1;
			10'b1101000000: counter[42] <= counter[42] + 1;
			10'b1101000001: counter[42] <= counter[42] + 1;
			10'b1101000010: counter[42] <= counter[42] + 1;
			10'b1101000011: counter[42] <= counter[42] + 1;
			10'b1101000100: counter[42] <= counter[42] + 1;
			10'b1101000101: counter[42] <= counter[42] + 1;
			10'b1101000110: counter[42] <= counter[42] + 1;
			10'b1101000111: counter[42] <= counter[42] + 1;
			10'b1101001000: counter[42] <= counter[42] + 1;
			10'b1101001001: counter[43] <= counter[43] + 1;
			10'b1101001010: counter[43] <= counter[43] + 1;
			10'b1101001011: counter[43] <= counter[43] + 1;
			10'b1101001100: counter[43] <= counter[43] + 1;
			10'b1101001101: counter[43] <= counter[43] + 1;
			10'b1101001110: counter[43] <= counter[43] + 1;
			10'b1101001111: counter[43] <= counter[43] + 1;
			10'b1101010000: counter[43] <= counter[43] + 1;
			10'b1101010001: counter[43] <= counter[43] + 1;
			10'b1101010010: counter[43] <= counter[43] + 1;
			10'b1101010011: counter[43] <= counter[43] + 1;
			10'b1101010100: counter[43] <= counter[43] + 1;
			10'b1101010101: counter[43] <= counter[43] + 1;
			10'b1101010110: counter[43] <= counter[43] + 1;
			10'b1101010111: counter[43] <= counter[43] + 1;
			10'b1101011000: counter[43] <= counter[43] + 1;
			10'b1101011001: counter[43] <= counter[43] + 1;
			10'b1101011010: counter[43] <= counter[43] + 1;
			10'b1101011011: counter[43] <= counter[43] + 1;
			10'b1101011100: counter[43] <= counter[43] + 1;
			10'b1101011101: counter[44] <= counter[44] + 1;
			10'b1101011110: counter[44] <= counter[44] + 1;
			10'b1101011111: counter[44] <= counter[44] + 1;
			10'b1101100000: counter[44] <= counter[44] + 1;
			10'b1101100001: counter[44] <= counter[44] + 1;
			10'b1101100010: counter[44] <= counter[44] + 1;
			10'b1101100011: counter[44] <= counter[44] + 1;
			10'b1101100100: counter[44] <= counter[44] + 1;
			10'b1101100101: counter[44] <= counter[44] + 1;
			10'b1101100110: counter[44] <= counter[44] + 1;
			10'b1101100111: counter[44] <= counter[44] + 1;
			10'b1101101000: counter[44] <= counter[44] + 1;
			10'b1101101001: counter[44] <= counter[44] + 1;
			10'b1101101010: counter[44] <= counter[44] + 1;
			10'b1101101011: counter[44] <= counter[44] + 1;
			10'b1101101100: counter[44] <= counter[44] + 1;
			10'b1101101101: counter[44] <= counter[44] + 1;
			10'b1101101110: counter[44] <= counter[44] + 1;
			10'b1101101111: counter[44] <= counter[44] + 1;
			10'b1101110000: counter[44] <= counter[44] + 1;
			10'b1101110001: counter[45] <= counter[45] + 1;
			10'b1101110010: counter[45] <= counter[45] + 1;
			10'b1101110011: counter[45] <= counter[45] + 1;
			10'b1101110100: counter[45] <= counter[45] + 1;
			10'b1101110101: counter[45] <= counter[45] + 1;
			10'b1101110110: counter[45] <= counter[45] + 1;
			10'b1101110111: counter[45] <= counter[45] + 1;
			10'b1101111000: counter[45] <= counter[45] + 1;
			10'b1101111001: counter[45] <= counter[45] + 1;
			10'b1101111010: counter[45] <= counter[45] + 1;
			10'b1101111011: counter[45] <= counter[45] + 1;
			10'b1101111100: counter[45] <= counter[45] + 1;
			10'b1101111101: counter[45] <= counter[45] + 1;
			10'b1101111110: counter[45] <= counter[45] + 1;
			10'b1101111111: counter[45] <= counter[45] + 1;
			10'b1110000000: counter[45] <= counter[45] + 1;
			10'b1110000001: counter[45] <= counter[45] + 1;
			10'b1110000010: counter[45] <= counter[45] + 1;
			10'b1110000011: counter[45] <= counter[45] + 1;
			10'b1110000100: counter[45] <= counter[45] + 1;
			10'b1110000101: counter[46] <= counter[46] + 1;
			10'b1110000110: counter[46] <= counter[46] + 1;
			10'b1110000111: counter[46] <= counter[46] + 1;
			10'b1110001000: counter[46] <= counter[46] + 1;
			10'b1110001001: counter[46] <= counter[46] + 1;
			10'b1110001010: counter[46] <= counter[46] + 1;
			10'b1110001011: counter[46] <= counter[46] + 1;
			10'b1110001100: counter[46] <= counter[46] + 1;
			10'b1110001101: counter[46] <= counter[46] + 1;
			10'b1110001110: counter[46] <= counter[46] + 1;
			10'b1110001111: counter[46] <= counter[46] + 1;
			10'b1110010000: counter[46] <= counter[46] + 1;
			10'b1110010001: counter[46] <= counter[46] + 1;
			10'b1110010010: counter[46] <= counter[46] + 1;
			10'b1110010011: counter[46] <= counter[46] + 1;
			10'b1110010100: counter[46] <= counter[46] + 1;
			10'b1110010101: counter[46] <= counter[46] + 1;
			10'b1110010110: counter[46] <= counter[46] + 1;
			10'b1110010111: counter[46] <= counter[46] + 1;
			10'b1110011000: counter[46] <= counter[46] + 1;
			10'b1110011001: counter[47] <= counter[47] + 1;
			10'b1110011010: counter[47] <= counter[47] + 1;
			10'b1110011011: counter[47] <= counter[47] + 1;
			10'b1110011100: counter[47] <= counter[47] + 1;
			10'b1110011101: counter[47] <= counter[47] + 1;
			10'b1110011110: counter[47] <= counter[47] + 1;
			10'b1110011111: counter[47] <= counter[47] + 1;
			10'b1110100000: counter[47] <= counter[47] + 1;
			10'b1110100001: counter[47] <= counter[47] + 1;
			10'b1110100010: counter[47] <= counter[47] + 1;
			10'b1110100011: counter[47] <= counter[47] + 1;
			10'b1110100100: counter[47] <= counter[47] + 1;
			10'b1110100101: counter[47] <= counter[47] + 1;
			10'b1110100110: counter[47] <= counter[47] + 1;
			10'b1110100111: counter[47] <= counter[47] + 1;
			10'b1110101000: counter[47] <= counter[47] + 1;
			10'b1110101001: counter[47] <= counter[47] + 1;
			10'b1110101010: counter[47] <= counter[47] + 1;
			10'b1110101011: counter[47] <= counter[47] + 1;
			10'b1110101100: counter[47] <= counter[47] + 1;
			10'b1110101101: counter[48] <= counter[48] + 1;
			10'b1110101110: counter[48] <= counter[48] + 1;
			10'b1110101111: counter[48] <= counter[48] + 1;
			10'b1110110000: counter[48] <= counter[48] + 1;
			10'b1110110001: counter[48] <= counter[48] + 1;
			10'b1110110010: counter[48] <= counter[48] + 1;
			10'b1110110011: counter[48] <= counter[48] + 1;
			10'b1110110100: counter[48] <= counter[48] + 1;
			10'b1110110101: counter[48] <= counter[48] + 1;
			10'b1110110110: counter[48] <= counter[48] + 1;
			10'b1110110111: counter[48] <= counter[48] + 1;
			10'b1110111000: counter[48] <= counter[48] + 1;
			10'b1110111001: counter[48] <= counter[48] + 1;
			10'b1110111010: counter[48] <= counter[48] + 1;
			10'b1110111011: counter[48] <= counter[48] + 1;
			10'b1110111100: counter[48] <= counter[48] + 1;
			10'b1110111101: counter[48] <= counter[48] + 1;
			10'b1110111110: counter[48] <= counter[48] + 1;
			10'b1110111111: counter[48] <= counter[48] + 1;
			10'b1111000000: counter[48] <= counter[48] + 1;
			10'b1111000001: counter[49] <= counter[49] + 1;
			10'b1111000010: counter[49] <= counter[49] + 1;
			10'b1111000011: counter[49] <= counter[49] + 1;
			10'b1111000100: counter[49] <= counter[49] + 1;
			10'b1111000101: counter[49] <= counter[49] + 1;
			10'b1111000110: counter[49] <= counter[49] + 1;
			10'b1111000111: counter[49] <= counter[49] + 1;
			10'b1111001000: counter[49] <= counter[49] + 1;
			10'b1111001001: counter[49] <= counter[49] + 1;
			10'b1111001010: counter[49] <= counter[49] + 1;
			10'b1111001011: counter[49] <= counter[49] + 1;
			10'b1111001100: counter[49] <= counter[49] + 1;
			10'b1111001101: counter[49] <= counter[49] + 1;
			10'b1111001110: counter[49] <= counter[49] + 1;
			10'b1111001111: counter[49] <= counter[49] + 1;
			10'b1111010000: counter[49] <= counter[49] + 1;
			10'b1111010001: counter[49] <= counter[49] + 1;
			10'b1111010010: counter[49] <= counter[49] + 1;
			10'b1111010011: counter[49] <= counter[49] + 1;
			10'b1111010100: counter[49] <= counter[49] + 1;
			10'b1111010101: counter[50] <= counter[50] + 1;
			10'b1111010110: counter[50] <= counter[50] + 1;
			10'b1111010111: counter[50] <= counter[50] + 1;
			10'b1111011000: counter[50] <= counter[50] + 1;
			10'b1111011001: counter[50] <= counter[50] + 1;
			10'b1111011010: counter[50] <= counter[50] + 1;
			10'b1111011011: counter[50] <= counter[50] + 1;
			10'b1111011100: counter[50] <= counter[50] + 1;
			10'b1111011101: counter[50] <= counter[50] + 1;
			10'b1111011110: counter[50] <= counter[50] + 1;
			10'b1111011111: counter[50] <= counter[50] + 1;
			10'b1111100000: counter[50] <= counter[50] + 1;
			10'b1111100001: counter[50] <= counter[50] + 1;
			10'b1111100010: counter[50] <= counter[50] + 1;
			10'b1111100011: counter[50] <= counter[50] + 1;
			10'b1111100100: counter[50] <= counter[50] + 1;
			10'b1111100101: counter[50] <= counter[50] + 1;
			10'b1111100110: counter[50] <= counter[50] + 1;
			10'b1111100111: counter[50] <= counter[50] + 1;
			10'b1111101000: counter[50] <= counter[50] + 1;
			10'b1111101001: counter[50] <= counter[50] + 1;
			10'b1111101010: counter[50] <= counter[50] + 1;
			10'b1111101011: counter[50] <= counter[50] + 1;
			10'b1111101100: counter[50] <= counter[50] + 1;
			10'b1111101101: counter[50] <= counter[50] + 1;
			10'b1111101110: counter[50] <= counter[50] + 1;
			10'b1111101111: counter[50] <= counter[50] + 1;
			10'b1111110000: counter[50] <= counter[50] + 1;
			10'b1111110001: counter[50] <= counter[50] + 1;
			10'b1111110010: counter[50] <= counter[50] + 1;
			10'b1111110011: counter[50] <= counter[50] + 1;
			10'b1111110100: counter[50] <= counter[50] + 1;
			10'b1111110101: counter[50] <= counter[50] + 1;
			10'b1111110110: counter[50] <= counter[50] + 1;
			10'b1111110111: counter[50] <= counter[50] + 1;
			10'b1111111000: counter[50] <= counter[50] + 1;
			10'b1111111001: counter[50] <= counter[50] + 1;
			10'b1111111010: counter[50] <= counter[50] + 1;
			10'b1111111011: counter[50] <= counter[50] + 1;
			10'b1111111100: counter[50] <= counter[50] + 1;
			10'b1111111101: counter[50] <= counter[50] + 1;
			10'b1111111110: counter[50] <= counter[50] + 1;
			10'b1111111111: counter[50] <= counter[50] + 1;
			default: a <= a ;
		endcase
		a <= 10'b0000000000; end
	else if (!signal & a!=10'b1111111111) begin
		a <= a + 1; end
	else if (!signal & a==10'b1111111111) begin
		a <= 10'b0000000000; end
	case(switch)
		6'b000001: ld = counter[1] ;
		6'b000010: ld = counter[2] ;
		6'b000011: ld = counter[3] ;
		6'b000100: ld = counter[4] ;
		6'b000101: ld = counter[5] ;
		6'b000110: ld = counter[6] ;
		6'b000111: ld = counter[7] ;
		6'b001000: ld = counter[8] ;
		6'b001001: ld = counter[9] ;
		6'b001010: ld = counter[10] ;
		6'b001011: ld = counter[11] ;
		6'b001100: ld = counter[12] ;
		6'b001101: ld = counter[13] ;
		6'b001110: ld = counter[14] ;
		6'b001111: ld = counter[15] ;
		6'b010000: ld = counter[16] ;
		6'b010001: ld = counter[17] ;
		6'b010010: ld = counter[18] ;
		6'b010011: ld = counter[19] ;
		6'b010100: ld = counter[20] ;
		6'b010101: ld = counter[21] ;
		6'b010110: ld = counter[22] ;
		6'b010111: ld = counter[23] ;
		6'b011000: ld = counter[24] ;
		6'b011001: ld = counter[25] ;
		6'b011010: ld = counter[26] ;
		6'b011011: ld = counter[27] ;
		6'b011100: ld = counter[28] ;
		6'b011101: ld = counter[29] ;
		6'b011110: ld = counter[30] ;
		6'b011111: ld = counter[31] ;
		6'b100000: ld = counter[32] ;
		6'b100001: ld = counter[33] ;
		6'b100010: ld = counter[34] ;
		6'b100011: ld = counter[35] ;
		6'b100100: ld = counter[36] ;
		6'b100101: ld = counter[37] ;
		6'b100110: ld = counter[38] ;
		6'b100111: ld = counter[39] ;
		6'b101000: ld = counter[40] ;
		6'b101001: ld = counter[41] ;
		6'b101010: ld = counter[42] ;
		6'b101011: ld = counter[43] ;
		6'b101100: ld = counter[44] ;
		6'b101101: ld = counter[45] ;
		6'b101110: ld = counter[46] ;
		6'b101111: ld = counter[47] ;
		6'b110000: ld = counter[48] ;
		6'b110001: ld = counter[49] ;
		6'b110010: ld = counter[50] ;
		default: ld = 8'b00000000; // Default case
	endcase
	end
end

assign led = ld;
assign gpio = ld2;
assign gpiob = y;
assign count = counter[0];

endmodule